library verilog;
use verilog.vl_types.all;
entity likeALU_tb is
end likeALU_tb;
